`include "fifo_common.sv"
`include "asynch_fifo.v"
`include "wr_tx.sv"
`include "wr_gen.sv"
`include "fifo_intrf.sv"
`include "wr_bfm.sv"
`include "wr_mon.sv"
`include "wr_cov.sv"
`include "wr_agent.sv"
`include "rd_tx.sv"
`include "rd_gen.sv"
`include "rd_bfm.sv"
`include "rd_mon.sv"
`include "rd_cov.sv"
`include "rd_agent.sv"
`include "fifo_sbd.sv"
`include "fifo_env.sv"
`include "fifo_assert.sv"
`include "top.sv"
